library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;

entity fulladder is
  port (
    x       : in  std_logic;
    y       : in  std_logic;
    c       : in  std_logic;
    z       : out std_logic;
    cout    : out std_logic
  );
end fulladder;

architecture structural_FA of fulladder is
signal xor0 : std_logic;
signal and0 : std_logic;
signal and1 : std_logic;
begin
  xor0_map  : xor_gate port map (x => x, y => y, z => xor0);
  xor1_map  : xor_gate port map (x => xor0, y => c, z => z);
  and0_map  : and_gate port map (x => x, y => y, z => and0);
  and1_map  : and_gate port map (x => xor0, y => c, z => and1);
  or0_map   : or_gate port map (x => and0, y => and1, z => cout);
end architecture structural_FA;

library ieee;
use ieee.std_logic_1164.all;

entity adder is
  port (
    A     : in std_logic_vector (31 downto 0);
    B     : in std_logic_vector (31 downto 0);
    R     : out std_logic_vector (31 downto 0)
  );
end adder;

architecture structural_adder of adder is
component fulladder
  port (
    x       : in  std_logic;
    y       : in  std_logic;
    c       : in  std_logic;
    z       : out std_logic;
    cout    : out std_logic
  );
end component fulladder;
signal C    : std_logic_vector (31 downto 0);
begin
  unit_first  : fulladder port map (x => A(0), y => B(0), c => '0', z => R(0), cout => C(0));
  unit_others : for i in 1 to 31 generate
  begin
    unit_map  : fulladder port map (x => A(i), y => B(i), c => C(i-1), z => R(i), cout => C(i));
  end generate unit_others;
end architecture structural_adder;
